`include "lib/defines.vh"
module EX(
    input wire clk,
    input wire rst,
    // input wire flush,
    input wire [`StallBus-1:0] stall,

    input wire [`ID_TO_EX_WD-1:0] id_to_ex_bus,

    output wire [`EX_TO_MEM_WD-1:0] ex_to_mem_bus,

    output wire data_sram_en,
    output wire [3:0] data_sram_wen,
    output wire [31:0] data_sram_addr,
    output wire [31:0] data_sram_wdata,
    output wire [`EX_TO_RF_BUS-1:0] ex_to_rf_bus,//Siri
    ///
    input wire [32:0] delay_ex
    ///
);

    reg [`ID_TO_EX_WD-1:0] id_to_ex_bus_r;
    reg [32:0] delay_ex_r;
    always @ (posedge clk) begin
        if (rst) begin
            id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
            delay_ex_r <=33'b0;
        end
        // else if (flush) begin
        //     id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
        // end
        else if (stall[2]==`Stop && stall[3]==`NoStop) begin
            id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
            delay_ex_r <=33'b0;
        end
        else if (stall[2]==`NoStop) begin
            id_to_ex_bus_r <= id_to_ex_bus;
            delay_ex_r<=delay_ex;
        end
    end

    wire [31:0] ex_pc, inst;
    wire [11:0] alu_op;
    wire [2:0] sel_alu_src1;
    wire [3:0] sel_alu_src2;
    // wire data_sram_en;         //
    // wire [3:0] data_sram_wen;  //
    wire rf_we;
    wire [4:0] rf_waddr;
    wire sel_rf_res;
    wire [31:0] rf_rdata1, rf_rdata2;
    //reg is_in_delayslot;

    assign {
        ex_pc,          // 148:117
        inst,           // 116:85
        alu_op,         // 84:83
        sel_alu_src1,   // 82:80
        sel_alu_src2,   // 79:76
        data_sram_en,    // 75
        data_sram_wen,   // 74:71
        rf_we,          // 70
        rf_waddr,       // 69:65
        sel_rf_res,     // 64
        rf_rdata1,         // 63:32
        rf_rdata2          // 31:0
    } = id_to_ex_bus_r;

    wire [31:0] imm_sign_extend, imm_zero_extend, sa_zero_extend;
    assign imm_sign_extend = {{16{inst[15]}},inst[15:0]};
    assign imm_zero_extend = {16'b0, inst[15:0]};
    assign sa_zero_extend = {27'b0,inst[10:6]};

    wire [31:0] alu_src1, alu_src2;
    wire [31:0] alu_result, ex_result;

    assign alu_src1 = sel_alu_src1[1] ? ex_pc :
                      sel_alu_src1[2] ? sa_zero_extend : rf_rdata1;

    assign alu_src2 = sel_alu_src2[1] ? imm_sign_extend :
                      sel_alu_src2[2] ? 32'h8 :
                      sel_alu_src2[3] ? imm_zero_extend : rf_rdata2;
    
    alu u_alu(
    	.alu_control (alu_op ),
        .alu_src1    (alu_src1    ),
        .alu_src2    (alu_src2    ),
        .alu_result  (alu_result  )
    );
    ////
    wire is_delay_slot_i;
    wire [31:0] link_address_o;  ///*****************************
   
    // wire [5:0]ld_and_st_op;
    assign 
    { 
    is_delay_slot_i,
    link_address_o
    }=delay_ex_r;
    
    wire [5:0] lw_sw_op; //lw_sw的前六位指令
    assign lw_sw_op=data_sram_en? inst[31:26]:6'b000000;
    assign data_sram_addr=data_sram_en? rf_rdata1+{{16{inst[15]}},inst[15:0]}:32'b0;
    assign data_sram_wdata=data_sram_en?rf_rdata2:32'b0;
    assign ex_result =is_delay_slot_i ? link_address_o:data_sram_en?data_sram_wdata:alu_result;
    ////
    
    // assign ex_result = (alu_op===12'b0)?alu_src1: data_sram_en? data_sram_wdata : alu_result;

     assign ex_to_mem_bus = {
        ex_pc,          // 81:50
        data_sram_en,    // 49
        data_sram_wen,   // 48:45
        sel_rf_res,     // 44
        rf_we,          // 43
        rf_waddr,       // 42:38
        lw_sw_op,   // 37:32
        ex_result       // 31:0
    };

    //Siri
    wire ex_to_rf_we;
    wire [4:0] ex_to_rf_waddr;
    wire [31:0] ex_to_rf_wdata;
    assign ex_to_rf_we =rf_we;
    assign ex_to_rf_waddr=rf_waddr;
    assign ex_to_rf_wdata=ex_result;
    assign ex_to_rf_bus={
        ex_to_rf_we,
        ex_to_rf_waddr,
        lw_sw_op,
        ex_to_rf_wdata
    };
    //Siri

    
    
endmodule